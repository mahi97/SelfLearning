entity datapath is
  port (
	clk, register_shift, register_load : in std_logic;
	register_out : out std_logic;
	register_in : in std_logic
  ) ;
end entity ; -- datapath

architecture rtl of datapath is

begin



end architecture ; -- rtl